module dependency_ctrl (
    
)