import rv32_pkg::*
module 